# ====================================================================
#
#      bootls.cdl
#
#      �ɶ���Ƽ������޹�˾��Ʒ�Ĳ�Ʒ��ʼ����ά�����ߡ�
#

cdl_package CYGPKG_BTOOLS {
    display		"BTOOLS Ӧ��"
	include_dir btools

	compile -library=libextras.a 	btools.c

	description "��Ʒ����ά������"

	make -priority 320 {
		<PREFIX>/bin/btools.elf : $(PREFIX)/lib/target.ld $(PREFIX)/lib/libtarget.a $(PREFIX)/lib/libextras.a
			@sh -c "mkdir -p $(dir $@)"
			$(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@
			$(COMMAND_PREFIX)strip $@ -o $(PREFIX)/bin/mini-btools.elf
	}

    cdl_option	CYGPKG_BTOOLS_AUTOEXEC {
        display		"�������Զ������ļ�ϵͳ��ִ��"
	    flavor        bool
        default_value 0
        description "�������Զ������ļ�ϵͳ��ִ��"
	}

    cdl_option	CYGPKG_BTOOLS_AUTO_INIT {
        display		"�������Զ���ɹ�����������"
	    flavor        bool
        default_value 0
        description "�������Զ���ɹ�����������"
	}
	
    cdl_component PRODUCE_BUILD_OPTIONS {
        display		"���ӵı���ѡ��"
        description "���ӵı���ѡ��"
		no_define
        flavor  none
        cdl_option PRODUCE_RADIUS_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package.
                These flags are used in addition
                to the set of global flags."
        }

        cdl_option PRODUCE_RADIUS_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }
    }

}
