# ====================================================================
#
#      hal_arm_at91sam9g20ek.cdl
#
#      ARM AT91SAM9G20-EK development board package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2006 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      danielh
# Contributors:
# Date:           2010-01-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_AT91SAM9G20EK {
    display       "Atmel AT91SAM9G20-EK board HAL"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_at91sam9g20ek.h
    include_dir   cyg/hal
    hardware
    description   "
	The AT91SAM9G20-EK HAL package provides the support needed to run
	eCos on an Atmel AT91SAM9G20-EK development board."

    compile       at91sam9g20ek_misc.c
    compile       at91sam9g20ek_mmu.c at91sam9g20ek_spi.c
    compile       -library=libextras.a at91sam9g20ek_flash.c at91sam9g20ek_redboot.c

    implements    CYGPKG_DEVS_FLASH_ATMEL_DATAFLASH_FLASH_DEV
    implements    CYGINT_HAL_ARM_ARCH_ARM9
    requires      { CYGHWR_HAL_ARM_AT91 == "AT91SAM9" }
    requires      { CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g20" }

    define_proc {
	puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_at91sam9g20ek.h>"
	puts $::cdl_header "/***** proc output start *****/"
	puts $::cdl_header "#include <pkgconf/hal_arm_at91sam9.h>"
	puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM926EJ-S\""
	puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Atmel AT91SAM9G20-EK\""
	puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
	puts $::cdl_header "/****** proc output end ******/"
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { (CYG_HAL_STARTUP == "RAM") ? \
		     "arm_at91sam9g20ek_ram" :
		     "arm_at91sam9g20ek_rom" }

	cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
	    display "Memory layout linker script fragment"
	    flavor data
	    no_define
	    define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
	    calculated { (CYGPKG_REDBOOT) ? \
		 "<pkgconf/mlt_arm_at91sam9g20ek_redboot.ldi>" :
		 "<pkgconf/mlt_arm_at91sam9g20ek_app.ldi>" }
	}

	cdl_option CYGHWR_MEMORY_LAYOUT_H {
	    display "Memory layout header file"
	    flavor data
	    no_define
	    define -file system.h CYGHWR_MEMORY_LAYOUT_H
	    calculated { (CYGPKG_REDBOOT) ? \
		 "<pkgconf/mlt_arm_at91sam9g20ek_redboot.h>" :
		 "<pkgconf/mlt_arm_at91sam9g20ek_app.h>" }
	}
    }
}
